-- André Luiz Rodrigues dos Santos RA1500759-UTFPR
-- Luí­s Henrique Beltã£o Santana RA906867-UTFPR
-- 20190411